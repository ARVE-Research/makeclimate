netcdf NAclimate {
dimensions:
	lon = 720 ;
	lat = 360 ;
	time = unlimited ;
variables:
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:actual_range = -180., 180. ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:actual_range = -90., 90. ;
	double time(time) ;
		time:avg_period = "0001-01-00 00:00:00" ;
		time:long_name = "time" ;
		time:actual_range = 0., 0. ;
		time:delta_t = "0000-01-00 00:00:00" ;
		time:standard_name = "time" ;
		time:coordinate_defines = "start" ;
		time:calendar = "proleptic_gregorian" ;
		time:note = "time coordinate refers to first day of month" ;
		time:units = "days since 1950-01-01 00:00:00" ;
		time:axis = "T" ;
	short elv(lat, lon) ;
		elv:long_name = "Elevation above mean sea level" ;
		elv:units = "m" ;
		elv:scale_factor = 1.f ;
		elv:add_offset = 0.f ;
		elv:_FillValue = -32768s ;
		elv:missing_value = -32768s ;
		elv:source = "ClimateNA v7.30" ;
		elv:actual_range = -196.f, 4893.f ;
		elv:_Storage = "chunked" ;
		elv:_ChunkSizes = 30, 30 ;
		elv:_DeflateLevel = 1 ;
	short tmp(time, lat, lon) ;
		tmp:long_name = "2m air temperature" ;
		tmp:units = "degC" ;
		tmp:scale_factor = 0.1f ;
		tmp:add_offset = 0.f ;
		tmp:_FillValue = -32768s ;
		tmp:missing_value = -32768s ;
		tmp:avg_period = "1950-2000" ;
		tmp:source = "ClimateNA v7.30" ;
		tmp:actual_range = -47.6f, 29.f ;
		tmp:_Storage = "chunked" ;
		tmp:_ChunkSizes = 360, 30, 30 ;
		tmp:_DeflateLevel = 1 ;
	short dtr(time, lat, lon) ;
		dtr:long_name = "Diurnal temperature range" ;
		dtr:units = "degC" ;
		dtr:scale_factor = 0.1f ;
		dtr:add_offset = 0.f ;
		dtr:_FillValue = -32768s ;
		dtr:missing_value = -32768s ;
		dtr:avg_period = "1950-2000" ;
		dtr:source = "ClimateNA v7.30" ;
		dtr:actual_range = -42.8f, 46.5f ;
		dtr:_Storage = "chunked" ;
		dtr:_ChunkSizes = 360, 30, 30 ;
		dtr:_DeflateLevel = 1 ;
	short pre(time, lat, lon) ;
		pre:long_name = "Total precipitation" ;
		pre:units = "mm" ;
		pre:scale_factor = 1.f ;
		pre:add_offset = 32767.f ;
		pre:_FillValue = -32768s ;
		pre:missing_value = -32768s ;
		pre:avg_period = "1950-2000" ;
		pre:source = "ClimateNA v7.30" ;
		pre:actual_range = 0.f, 1840.f ;
		pre:_Storage = "chunked" ;
		pre:_ChunkSizes = 360, 30, 30 ;
		pre:_DeflateLevel = 1 ;
	short wet(time, lat, lon) ;
		wet:long_name = "Fraction of days in the month with > 0.1mm precipitation" ;
		wet:units = "fraction" ;
		wet:scale_factor = 0.01f ;
		wet:add_offset = 0.f ;
		wet:_FillValue = -32768s ;
		wet:missing_value = -32768s ;
		wet:avg_period = "1950-2000" ;
		wet:source = "modeled on climateNA v7.30 precip using CRU TS4.06 empirical relationship" ;
		wet:actual_range = 0.f, 1.f ;
		wet:_Storage = "chunked" ;
		wet:_ChunkSizes = 360, 30, 30 ;
		wet:_DeflateLevel = 1 ;
	short cld(time, lat, lon) ;
		cld:long_name = "Total cloud cover fraction" ;
		cld:units = "fraction" ;
		cld:scale_factor = 0.1f ;
		cld:add_offset = 0.f ;
		cld:_FillValue = -32768s ;
		cld:missing_value = -32768s ;
		cld:avg_period = "1950-2000" ;
		cld:source = "CHELSA v2.1" ;
		cld:actual_range = 4.5f, 90.7f ;
		cld:_Storage = "chunked" ;
		cld:_ChunkSizes = 360, 30, 30 ;
		cld:_DeflateLevel = 1 ;
	short wnd(time, lat, lon) ;
		wnd:long_name = "10m windspeed" ;
		wnd:units = "m s-1" ;
		wnd:scale_factor = 0.001f ;
		wnd:add_offset = 0.f ;
		wnd:_FillValue = -32768s ;
		wnd:missing_value = -32768s ;
		wnd:avg_period = "1950-2000" ;
		wnd:source = "CHELSA v2.1" ;
		wnd:actual_range = 0.284f, 22.082f ;
		wnd:_Storage = "chunked" ;
		wnd:_ChunkSizes = 360, 30, 30 ;
		wnd:_DeflateLevel = 1 ;
	short lght(time, lat, lon) ;
		lght:long_name = "Lightning stroke density" ;
		lght:units = "km-2 d-1" ;
		lght:scale_factor = 1.e-05f ;
		lght:add_offset = 0.32767f ;
		lght:_FillValue = -32768s ;
		lght:missing_value = -32768s ;
		lght:avg_period = "2012-2021" ;
		lght:source = "WGLC" ;
		lght:actual_range = 2.980232e-08f, 0.39123f ;
		lght:_Storage = "chunked" ;
		lght:_ChunkSizes = 360, 30, 30 ;
		lght:_DeflateLevel = 1 ;

// global attributes:
		:Conventions = "COARDS, CF-1.11" ;
		:title = "ANOMTYPE global climate, 30m grid" ;
		:note = "based on ClimateNA v7.30, CHELSA 2.1, and WGLC with anomalies from ModelE-LM" ;
		:node_offset = 1 ;
}
