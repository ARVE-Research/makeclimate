netcdf NAclimate {
dimensions:
	x = 1539 ;
	y = 1533 ;
	time = unlimited ;
variables:
	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:units = "meter" ;
		x:axis = "X" ;
		x:actual_range = -4350000., 3345000. ;
	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:units = "meter" ;
		y:axis = "Y" ;
		y:actual_range = -3885000., 3780000. ;
	double time(time) ;
		time:avg_period = "0001-01-00 00:00:00" ;
		time:long_name = "time" ;
		time:actual_range = 0., 0. ;
		time:delta_t = "0000-01-00 00:00:00" ;
		time:standard_name = "time" ;
		time:coordinate_defines = "start" ;
		time:calendar = "proleptic_gregorian" ;
		time:note = "time coordinate refers to first day of month" ;
		time:units = "days since 1836-01-01 00:00:00" ;
		time:axis = "T" ;
	double lon(y, x) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:actual_range = -179.999908447266, 179.99967956543 ;
		lon:grid_mapping = "crs" ;
		lon:_Storage = "chunked" ;
		lon:_ChunkSizes = 25, 25 ;
		lon:_DeflateLevel = 1 ;
	double lat(y, x) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:actual_range = 5.48972606658936, 84.4052429199219 ;
		lat:grid_mapping = "crs" ;
		lat:_Storage = "chunked" ;
		lat:_ChunkSizes = 25, 25 ;
		lat:_DeflateLevel = 1 ;
	short elv(y, x) ;
		elv:long_name = "Elevation above mean sea level" ;
		elv:units = "m" ;
		elv:scale_factor = 1.f ;
		elv:add_offset = 0.f ;
		elv:_FillValue = -32768s ;
		elv:missing_value = -32768s ;
		elv:source = "ClimateNA v7.30" ;
		elv:actual_range = -196.f, 4893.f ;
		elv:grid_mapping = "crs" ;
		elv:_Storage = "chunked" ;
		elv:_ChunkSizes = 25, 25 ;
		elv:_DeflateLevel = 1 ;
	short tmp(time, y, x) ;
		tmp:long_name = "2m air temperature" ;
		tmp:units = "degC" ;
		tmp:scale_factor = 0.1f ;
		tmp:add_offset = 0.f ;
		tmp:_FillValue = -32768s ;
		tmp:missing_value = -32768s ;
		tmp:avg_period = "1950-2000" ;
		tmp:source = "ClimateNA v7.30" ;
		tmp:actual_range = -47.6f, 29.f ;
		tmp:grid_mapping = "crs" ;
		tmp:_Storage = "chunked" ;
		tmp:_ChunkSizes = 360, 25, 25 ;
		tmp:_DeflateLevel = 1 ;
	short dtr(time, y, x) ;
		dtr:long_name = "Diurnal temperature range" ;
		dtr:units = "degC" ;
		dtr:scale_factor = 0.1f ;
		dtr:add_offset = 0.f ;
		dtr:_FillValue = -32768s ;
		dtr:missing_value = -32768s ;
		dtr:avg_period = "1950-2000" ;
		dtr:source = "ClimateNA v7.30" ;
		dtr:actual_range = -42.8f, 46.5f ;
		dtr:grid_mapping = "crs" ;
		dtr:_Storage = "chunked" ;
		dtr:_ChunkSizes = 360, 25, 25 ;
		dtr:_DeflateLevel = 1 ;
	short pre(time, y, x) ;
		pre:long_name = "Total precipitation" ;
		pre:units = "mm" ;
		pre:scale_factor = 1.f ;
		pre:add_offset = 32767.f ;
		pre:_FillValue = -32768s ;
		pre:missing_value = -32768s ;
		pre:avg_period = "1950-2000" ;
		pre:source = "ClimateNA v7.30" ;
		pre:actual_range = 0.f, 1840.f ;
		pre:grid_mapping = "crs" ;
		pre:_Storage = "chunked" ;
		pre:_ChunkSizes = 360, 25, 25 ;
		pre:_DeflateLevel = 1 ;
	short wet(time, y, x) ;
		wet:long_name = "Fraction of days in the month with > 0.1mm precipitation" ;
		wet:units = "fraction" ;
		wet:scale_factor = 0.01f ;
		wet:add_offset = 0.f ;
		wet:_FillValue = -32768s ;
		wet:missing_value = -32768s ;
		wet:avg_period = "1950-2000" ;
		wet:source = "modeled on climateNA v7.30 precip using CRU TS4.06 empirical relationship" ;
		wet:actual_range = 0.f, 1.f ;
		wet:grid_mapping = "crs" ;
		wet:_Storage = "chunked" ;
		wet:_ChunkSizes = 360, 25, 25 ;
		wet:_DeflateLevel = 1 ;
	short cld(time, y, x) ;
		cld:long_name = "Total cloud cover fraction" ;
		cld:units = "fraction" ;
		cld:scale_factor = 0.1f ;
		cld:add_offset = 0.f ;
		cld:_FillValue = -32768s ;
		cld:missing_value = -32768s ;
		cld:avg_period = "1950-2000" ;
		cld:source = "CHELSA v2.1" ;
		cld:actual_range = 4.5f, 90.7f ;
		cld:grid_mapping = "crs" ;
		cld:_Storage = "chunked" ;
		cld:_ChunkSizes = 360, 25, 25 ;
		cld:_DeflateLevel = 1 ;
	short wnd(time, y, x) ;
		wnd:long_name = "10m windspeed" ;
		wnd:units = "m s-1" ;
		wnd:scale_factor = 0.001f ;
		wnd:add_offset = 0.f ;
		wnd:_FillValue = -32768s ;
		wnd:missing_value = -32768s ;
		wnd:avg_period = "1950-2000" ;
		wnd:source = "CHELSA v2.1" ;
		wnd:actual_range = 0.284f, 22.082f ;
		wnd:grid_mapping = "crs" ;
		wnd:_Storage = "chunked" ;
		wnd:_ChunkSizes = 360, 25, 25 ;
		wnd:_DeflateLevel = 1 ;
	short lght(time, y, x) ;
		lght:long_name = "Lightning stroke density" ;
		lght:units = "km-2 d-1" ;
		lght:scale_factor = 1.e-05f ;
		lght:add_offset = 0.32767f ;
		lght:_FillValue = -32768s ;
		lght:missing_value = -32768s ;
		lght:avg_period = "2012-2021" ;
		lght:source = "WGLC" ;
		lght:actual_range = 2.980232e-08f, 0.39123f ;
		lght:grid_mapping = "crs" ;
		lght:_Storage = "chunked" ;
		lght:_ChunkSizes = 360, 25, 25 ;
		lght:_DeflateLevel = 1 ;
	char lambert_azimuthal_equal_area ;
		lambert_azimuthal_equal_area:grid_mapping_name = "lambert_azimuthal_equal_area" ;
		lambert_azimuthal_equal_area:false_easting = 0. ;
		lambert_azimuthal_equal_area:false_northing = 0. ;
		lambert_azimuthal_equal_area:latitude_of_projection_origin = 50. ;
		lambert_azimuthal_equal_area:longitude_of_projection_origin = -100. ;
		lambert_azimuthal_equal_area:long_name = "CRS definition" ;
		lambert_azimuthal_equal_area:longitude_of_prime_meridian = 0. ;
		lambert_azimuthal_equal_area:semi_major_axis = 6378137. ;
		lambert_azimuthal_equal_area:inverse_flattening = 298.257223563 ;
		lambert_azimuthal_equal_area:spatial_ref = "PROJCS[\"North_America_Lambert_Azimuthal_Equal_Area\",GEOGCS[\"WGS 84\",DATUM[\"WGS_1984\",SPHEROID[\"WGS 84\",6378137,298.257223563],AUTHORITY[\"EPSG\",\"6326\"]],PRIMEM[\"Greenwich\",0,AUTHORITY[\"EPSG\",\"8901\"]],UNIT[\"degree\",0.0174532925199433]],PROJECTION[\"Lambert_Azimuthal_Equal_Area\"],PARAMETER[\"latitude_of_center\",50],PARAMETER[\"longitude_of_center\",-100],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]],AXIS[\"Easting\",EAST],AXIS[\"Northing\",NORTH]]" ;
		lambert_azimuthal_equal_area:GeoTransform = "-4350000 5000 0 3780000 0 -5000 " ;
	int crs ;
		crs:grid_mapping_name = "lambert_azimuthal_equal_area" ;
		crs:proj_params = "+proj=laea +lat_0=50 +lon_0=-100 +x_0=0 +y_0=0 +datum=WGS84 +units=m +no_defs" ;

// global attributes:
		:Conventions = "COARDS, CF-1.11" ;
		:title = "ANOMTYPE climate for North America, 5km LAEA grid, v. 1.0" ;
		:note = "based on ClimateNA v7.30, CHELSA 2.1, WGLC, and 20th Century Reanalysis" ;
		:node_offset = 1 ;
}
